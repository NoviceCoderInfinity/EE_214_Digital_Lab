library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity students is
	port( inp:in std_logic_vector(4 downto 0);
		reset,clock:in std_logic;
		outp: out std_logic);
end students;

architecture bhv of students is

type state is (rst,s1,s2,s3,s4,s5,s6,s7); 
signal y_present,y_next: state:=rst;

begin
clock_proc:process(clock,reset)
begin
	if(clock='1' and clock' event) then
		if(reset='1') then
			y_present<= rst; 
		else
			y_present<= y_next;
		end if;
	end if;
	
end process;
state_transition_proc:process(inp,y_present)
begin
	case y_present is
		when rst=>
			if(unsigned(inp)=19) then 
				y_next<= s1;
			else
				y_next<= rst;
			end if;
		when s1=>
			if(unsigned(inp)=20) then 
				y_next<= s2;
			else
				y_next<= s1;
			end if;
		when s2=>
			if(unsigned(inp)=21) then 
				y_next<= s3;
			else
				y_next<= s2;
			end if;
		when s3=>
			if(unsigned(inp)=4) then 
				y_next<= s4;
			else
				y_next<= s3;
			end if;
		when s4=>
			if(unsigned(inp)=5) then 
				y_next<= s5;
			else
				y_next<= s4;
			end if;
		when s5=>
			if(unsigned(inp)=14) then 
				y_next<= s6;
			else
				y_next<= s5;
			end if;
		when s6=>
			if(unsigned(inp)=20) then 
				y_next<= s7;
			else
				y_next<= s6;
			end if;
		when s7=>
			if(unsigned(inp)=19) then 
				y_next<= s1;
			else
				y_next<= s7;
			end if;
	end case;
end process;

output_proc: process(y_present, y_next)
begin
	case y_present is
		when rst=>
			outp <= '0';
		when s1=>
			outp <= '0';
		when s2=>
			outp <= '0';
		when s3=>
			outp <= '0';
		when s4=>
			outp <= '0';
		when s5=>
			outp <= '0';
		when s6=>
			outp <= '0';
		when s7=>
			if(y_next = s7) then
				outp <= '0';
			else
				outp <= '1';
			end if;
	end case;
end process;
end bhv;